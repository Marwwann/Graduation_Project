.param Len=1e-06
.param sb=1.0